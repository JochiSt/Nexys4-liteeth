../modules/Ethernet/build/gateware/liteeth_core.vhdl
../../modules/Ethernet/liteeth/liteeth_core.vhdl
../../modules/Ethernet/liteeth/build/gateware/liteeth_core.vhdl